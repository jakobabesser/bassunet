BZh91AY&SY���� �߀Px����������`_|����8׃�
� 6�C@w���aT��	@	�JyS�'����`��i���=U*��`�M44�d�4�ɦ��0&&�	�&L�&	�����@T�� `     �$#Jz�(��2 @�i��Ddh�O�yS��M����f)�^����
(�9��R�:7|���I!]ꢐ*'��M�ar��\X!��8�HAUL��H{ӿ���J���^^�4��
��e���?k@�������ʞ��&S�~������f��A�<N,�0��$�6�m�l�\��E�tR�B@�fI����-2�B7m�Z6�)%���A2�0��$mn�)�H�!���Di	5!(�).BZ��&;'���f�4ZI��cT������$>8l�s'"�s���Mg��WAU<O)�<���Qq�����U�X��$���ыq76` $݀n͋��Ȳɶ��n�۫@BHH0 r��b��ZҀ��"�I�- ���B� 0� ����-�� /N��V?b��!�O�e�����x(0�w�݊�ஊ&�H��j�2 �����E"@��ц�<�`��9���a�w��!\����9o���N3lbSRYkY�͖Kv��0��fw%��˟>sf�	��Vm�����"�B�*�!8V����Dڑ�B�r	�B�� x[+L<q#�N�!�� OF���ׂ�L|O+}4�K��Lq3�t�奀LՂDVQ��t�	G�D1U�Ӕҧ��=$��iS|p�s75u3S�
M����Q|�db���i��w7e�p���[&��zwe\�9�+9�ؖ�sF�#Rm+^�9bo�Silq�Z�Ц�JY!��!ѹɾ�$2�E��7m��-�քCD34+��!�A@))�V�(Vg֌h���H�1�զ��B���Ɲ"��\��i�`L�fαi����v�F�"�L�ѹ���Jp!��&a�i�Lb�}�&�oŀ'��JCC��#��jK��x&��a��L�i6ӆF�53�Fu�B�G�d��J^� (���g볦��Q�;zbs�n������H߇k��ت���5�t��Hۘ��$�f���%\l���iYf]�]���<�#{+���H6��iV�� � ��ccO#�Gz@�1,m��m�U�m�H� ^3����[k���EΊGQ�C;�5dA�0�m���i"Vj�=`�'EVq߀��0[�ھp���8��3I�[����^��JCC+DD*�·me�+c��(T�MN""��B����E���S��*�C�&s:�]E��ġ�7�����;�<f�4��*�;!k����g!��D��ԭ.�o"���8c%w%J�uD�EM��d���6�j�Q��I��.YÎ&۬��v\̓_� O+�ڠ�qq��P�!I�DM���;��m1{�*�/���il��z���TT����EVvu���j�-XV�Q���+{��"�qL��
��A0TVZҹd��k
�+�9̙��WM��n�'u�����n��|N���!��x�)Q�2aVFӨ�gy���[��Q��LT6�K�$��gx ����6�ul�F���P��f�hv�xx*��V3H��D�x*��3y�l�Y��ghX�d�{̮�挀W')�bDsaoi��ͧvwXx��ؽ�{��9���]%U[0W�=�^�5���p�w^ 0�k���eq�C������[�˵l�"Whv�{Ձ�J�eؾg-��ђ&��|�M'?�z�����I	$� (��TS���*��Ol*ՀQ�aaUTEQVHTAURkTTX#�LE��o�y`������0�@ja���"c�Ҳ��^���YM����2�ł����(s��Q�e�BQ,EC
Y�#h*�AGTfe	��z�YnC-��D]Q����@P�U� j������3�|�_��'�	O�?������?��������{a)�1Jx��:9�?�h=��k"�Ƹ/���8b�]]S��rcR�E2C�23p�ܾ��x��7����$B�Jm}D>��n��p`C��d?6ߖ�p����aݰ�TOC��UӒ����������OX/y� ������y�o��(��e�܂IXa�N���v&=��-J�Z���^}�pc��PP�@��B(�D�*�BB��e�,"���Ab`H�D�Ŋ$H"b)2����CL�ef@�6/W���AcQ�m��m�Z����D���21�s�ǈg������gM�����<Cc��Bkǎ l?M���Ә��\� T�XRz��<�Տ�z�S�=�˦aв�d�=����t��&�����ǫ��w��������&��9�?e��_3�f���Q� ��^@F�y�TS�l|jE�����j^���X�-��3��B�m����V�!�[K�s,�.� �,X9yfpn.)��Y�vY�� !���b.+�]ȏs�A�#����5j��� k<<�@�ܓ�;UE<}�� ��<x����q��f���
���<����C�SF��+�,t�>>o���Mw T�B�"y ��>��<E9"n��>&^MF�a�AېbrS"G`Q�����),B��6=��V�p��ݴvgd3����߰.�c�b�u5kԪ)���r��E�[[��}�������ǡ���* B���"{_ m��{D�
�F'�g�� ̂�=�8���9ۥ(]�:8��La����91�8B,��Vа=�1���=?!w$S�		
L�